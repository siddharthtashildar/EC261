module nor_not(input a, output y);
    nor (y, a, a);
endmodule
