`timescale 1ns/1ps

module tb_mux_testrun;

    reg I0, I1, I2, I3, I4, I5, I6, I7;
    reg S0, S1, S2;
    wire output_wire;

    
    mux uut (
        .I0(I0), .I1(I1), .I2(I2), .I3(I3),
        .I4(I4), .I5(I5), .I6(I6), .I7(I7),
        .S0(S0), .S1(S1), .S2(S2),
        .output_wire(output_wire)
    );



    initial begin
        
        $dumpfile("wave.vcd");
        $dumpvars(0, tb_mux_testrun);
        
        I0 = 0; I1 = 1; I2 = 0; I3 = 1;
        I4 = 0; I5 = 1; I6 = 0; I7 = 1;

        $display("Time | S2 S1 S0 | Output | Selected Input");

        S2=0; S1=0; S0=0; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=0; S1=0; S0=1; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=0; S1=1; S0=0; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=0; S1=1; S0=1; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=1; S1=0; S0=0; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=1; S1=0; S0=1; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=1; S1=1; S0=0; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        S2=1; S1=1; S0=1; #10;
        $display("Selected: I0=%b I1=%b I2=%b I3=%b I4=%b I5=%b I6=%b I7=%b", 
                 (S2==0 && S1==0 && S0==0), (S2==0 && S1==0 && S0==1), (S2==0 && S1==1 && S0==0), (S2==0 && S1==1 && S0==1),
                 (S2==1 && S1==0 && S0==0), (S2==1 && S1==0 && S0==1), (S2==1 && S1==1 && S0==0), (S2==1 && S1==1 && S0==1));

        $finish;
    end


    initial begin
        $monitor("%4t |  %b  %b  %b  |   %b", 
                 $time, S2, S1, S0, output_wire);
    end

endmodule