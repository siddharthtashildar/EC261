
module ring_counter_4bit (
    input clk,
    input rst,
    output reg [3:0] q
);
    always @(posedge clk or posedge rst) begin
        if (rst)
            q <= 4'b1000;              // Start with only one '1'
        else
            q <= {q[2:0], q[3]};       // Rotate left
    end
endmodule
