module johnson_counter_4bit (
    input clk,
    input rst,
    output reg [3:0] q
);
    always @(posedge clk or posedge rst) begin
        if (rst)
            q <= 4'b0000;                // start with all zeros
        else
            q <= {~q[0], q[3:1]};        // twisted feedback
    end
endmodule
